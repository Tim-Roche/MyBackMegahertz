module computer();
endmodule